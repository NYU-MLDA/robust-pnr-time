/home/abc586/freepdk-45nm/rtk-tech.lef