/home/abc586/freepdk-45nm/stdcells.lef